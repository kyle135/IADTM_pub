///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
//
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`default_nettype none
module reset_synchronizer #(
	parameter int	DEPTH		= 3,
	parameter bit	POLARITY	= 1
)  (//--------------------------------------------------------------//-------------------------------------------------
	//																//
	//--------------------------------------------------------------//-------------------------------------------------
	input	wire	source_rst,										//
	//--------------------------------------------------------------//-------------------------------------------------
	//																//
	//--------------------------------------------------------------//-------------------------------------------------
	input	wire	target_clk,										//
	output	wire	target_rst										//
);
//
	reg	[DEPTH] shift_reg;
	
	always_ff @(posedge target_clk ) begin
		if ( source_rst == POLARITY )	shift_reg	<= { DEPTH { POLARITY } };
		else							shift_reg	<= { shift_reg[DEPTH-2:0], source_rst };
	end
	//

	assign target_rst  = shift_reg[DEPTH-1];

endmodule : reset_synchronizer
`default_nettype wire
