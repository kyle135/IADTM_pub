`ifndef DESIGN_VH
    `define DESIGN_VH


`include "design_functions.vh"



`endif
