




module ProcessorStatus(


);



    // R3000 (MIPS I) status register
    typedef union packed {
        logic [31:0] ProcessorStatus_w;
        struct packed {
            logic [1:0] B31_30;  // [31:30] Unused
            logic       CU1;     // [   29] Coprocessor I usable: 1 to use FPA if you have it, 0 to disable. When 0, all FPA instructions cause an exception. While it's obviously a bad idea to enable FPA instructions if your CPU lacks FPA hardware, it can be useful to turn off an FPA even when you haye one.
            logic       CU0;     // [   28] Coprocessor 0 usable: Set I to be able to use some nominally privileged instructions in user mode. You don't want to do this. The CPU control instructions encoded as coprocessor 0 type are always usable in kernel mode, regardless of the setting of this bit.
            logic [1:0] B27_26;  // [27:26] Unused
            logic       RE;      // [   25] Reverse endianness in user mode: The MIPS processors can be configured, at reset time, with either endianness. Since human beings are perverse, there are now two universes of MIPS implementation: DEC and Windows NT are little-endian; SGI and their UNIX world are big-endian. Embedded applications originally showed a strong big-endian bias but are now thoroughly mixed. It could be a useful feature in an operating system to be able to run software from the opposite universe; the RE bit makes it possible. When RE is active, user-privilege software runs as if the CPU had been configured with the opposite endianness.
            logic [1:0] B24_23;  // [24:23] Unused
            logic       BEV;     // [   22] Boot exception vectors: When BEV == I, the CPU uses the ROM (ksegl) space exception entry point. BEV is usually set to 0 in running systems.
            logic       TS;      // [   21] TLB shutdown: See Chapter 6 for details. TS gets set if a program address simultaneously matches two TLB entries, which is certainly a sign of something horribly wrong in the OS soft- ware. Prolonged operation in this state, in some implementa- tions, could cause internal contention and damage to some chips, so the TLB ceases to match anything. TLB shutdown is terminal and can be cleared only by a hardware reset. Some MIPS CPUs have foolproof TLB hardware and may not implement this bit. Ön IDT R3051 family CPUs you can inspect this bit following hardware reset, and it will be set if and only if the CPU lacks a TLB (the memory management hardware). This test is not reliable across all implementations.
            logic       PE;      // [   20] Set if a cache parity error has occurred. No exception is generated by this condition, which is really only useful for diagnostics. The MIPS architecture has cache diagnostic facilities because earlier versions of the CPU used external caches, and signal timing on the cache buses was at the limits of technology. For those implementations the cache parity error bit was an essential design debug tool.
            logic       CM;      // [   19] This shows the result of the last load operation performed with the D-cache isolated. CM is set if the cache really contained data for the addressed memory location (i.e., if the load would have hit in the cache even if the cache had not been isolated).
            logic       PZ;      // [   18] When set, cache parity bits are written as zero and not checked. This is a fossil from CPUs with external caches, where it allowed confident designers to dispense with the external memory that held the cache parity bits, saving a little money. You won't use this if the CPU has on-chip caches.
            //  Swap caches and isolate (data) cache: These are cache mode bits for cache management and diagnostics;
            logic       SwC;     // [   17] When SR(SMC) is set, the roles of the I-cache and the D-cache are reversed so that you can access and invalidate I-cache entries.
            logic       IsC;     // [   16] When SR(IsC) is set, all loads and stores access only the data cache and never memory; in this mode a partial-word store invalidates the cache entry. 
            logic [7:0] IM;      // [15: 8] Interrupt mask: An 8-bit field defining which interrupt sources, when active, will be allowed to cause an exception. Six of the interrupt sources are generated by signals from outside the CPU core (one may be used by the FPA, which although it lives on the same chip is logically external); the other two are the software-writable interrupt bits in the Cause register. The 32-bit CPUs with floating-point hardware use one of the CPU interruptsto signal floating-point exceptions; MIPS III and subsequent CPUs usually have an interval timer as part of the co- processor 0 features, and timer events are signalled on the high- est interrupt bit. Otherwise, interrupts are signalled from out- side the CPU chip. No interrupt prioritization is provided for you: The hardware treats all interrupt bits the same. See Section 5.8 for details.
            logic [1:0] B07_06;  // [ 7: 6] Unused
            logic       KUo;     // [    5] KU old. On an exception the KUp bit is saved
            logic       IEo;     // [    4] IE old. On an exception the IEP bit is saved
            // On an exception, the hardware takes the values ofKUc and IEC and saves them here at the same time as changing the values of KUc, IEc to [1, 0] (kernel mode, interrupts disabled). The instruction rfe can be used to copy KUp, IEP back into KUc, IEc.
            logic       KUp;     // [    3] KU previous
            logic       IEp;     // [    2] IE previous
            // These are the two basic CPU protection bits.            
            logic       KUc;     // [    1] KUC is set I when running with kernel privileges, 0 for user mode. In kernel mode you can get at the whole program address space and use privileged (coprocessor 0) instructions. In user mode you are restricted to program addresses between zero and 0x7FFF FFFF and can't run privileged instructions; attempts to break the rules result in an exception.
            logic       IEc;     // [    0] IEC is set 0 to prevent the CPU taking an interrupt, 1 to enable.
        } ProcessorStatus_s;
    } R3000_ProcessorStatus_t;


endmodule : ProcessorStatus