
module BehavioralAddRippleCarry
#(  //--------------------------------------//---------------------------------
    // Parameters                           // Description(s)
    //--------------------------------------//---------------------------------
    parameter int    N     = 32             //
)  (//--------------------------------------//---------------------------------
    // Inputs                               // Description(s)
    //--------------------------------------//---------------------------------
    input  wire [N-1:0] a,                  //
    input  wire [N-1:0] b,                  //
    input  wire         carry_in,           //
    //--------------------------------------//---------------------------------
    // Outputs                              // Description(s)
    //--------------------------------------//---------------------------------
    output reg  [N-1:0] c,                  //
    output reg          carry_out           //
);

    //-------------------------------------------------------------------------
    // Local Signals
    //-------------------------------------------------------------------------
    reg [N-1:0] carry;

    //-------------------------------------------------------------------------
    // Combinational Logic
    //-------------------------------------------------------------------------
    always@* c         = a ^ b ^ {carry[N-2:0], carry_in};
    always@* carry     = {carry[N-2:0], carry_in} & (a | b) | (a & b);
    always@* carry_out = carry[N-1];

endmodule : BehavioralAddRippleCarry
