//---------------------------------------------------------------------------------------
// Company: It's All Digital To Me
// Engineer: Kyle D. Gilsdorf
// Create Date: 09/21/2013
// Design Name: Structural Logical Less Than (by n-bits)
// Unit Name: Logical
// Module Name: StructuralLogicalGT
// Project Name: BasicCombinationalLogic
// Dependencies: None
//---------------------------------------------------------------------------------------
`default_nettype none
module StructuralLogicalLT
#(  //----------------------------------//-------------------------------------
    // Parameter(s)                     // Description(s)
    //----------------------------------//-------------------------------------
    parameter integer N = 8             // The number of bits of the operands.
)  (//----------------------------------//-------------------------------------
    // Input(s)                         // Description(s)
    //----------------------------------//-------------------------------------
    input  wire [N-1:0] a,              // Operand A
    input  wire [N-1:0] b,              // Operand B
    //----------------------------------//-------------------------------------
    // Output(s)                        // Description(s)
    //----------------------------------//-------------------------------------
    output reg           c               // Result C
);

    //-------------------------------------------------------------------------
    // Local Signals
    //-------------------------------------------------------------------------
    wire [N-1:0] an;
    wire [(N/4)-1:0] lt;
    wire [(N/4)-1:0] gt;
    wire [(N/4)-1:0] eq;
    //-------------------------------------------------------------------------
    // Combinational Logic
    //-------------------------------------------------------------------------

    //-------------------------------------------------------------------------
    // Module instance(s)
    //-------------------------------------------------------------------------

    genvar i;
    generate
    for (i = 0; i < (N/4); i = i + 1) begin : LT_BLOCK
        assign eq[i] = 
            ~(a[(i*4)+3] ^ b[(i*4)+3]) & 
            ~(a[(i*4)+2] ^ b[(i*4)+2]) &
            ~(a[(i*4)+1] ^ b[(i*4)+1]) &
            ~(a[(i*4)+0] ^ b[(i*4)+0]);
        //  Greater Than
        // .---.---.---.---.---.---.---.---.
        // | a | a | a | a | b | b | b | b |
        // | 3 | 2 | 1 | 0 | 3 | 2 | 1 | 0 |
        // :---+---+---+---+---+---+---+---:
        // | 1 | x | x | x | 0 | x | x | x | T
        // | 0 | 1 | x | x | 0 | 0 | x | x | T 
        // | 0 | 0 | 1 | x | 0 | 0 | 0 | x | T 
        // | 0 | 0 | 0 | 1 | 0 | 0 | 0 | 0 | T
        // '---'---'---'---'---'---'---'---'
        assign gt[i] =
            ( a[(i*4)+3] & a[(i*4)+2] & a[i+1] & a[(i*4)+0] & ~b[(i*4)+3] & ~b[(i*4)+2] & ~b[(i*4)+1] & ~b[(i*4)+0]) |
            ( a[(i*4)+3] & a[(i*4)+2] & a[i+1]              & ~b[(i*4)+3] & ~b[(i*4)+2] & ~b[(i*4)+1]) |
            ( a[(i*4)+3] & a[(i*4)+2]                       & ~b[(i*4)+3] & ~b[(i*4)+2]) |
            ( a[(i*4)+3]                                    & ~b[(i*4)+3]);

        //  Less Than
        // .---.---.---.---.---.---.---.---.
        // | a | a | a | a | b | b | b | b |
        // | 3 | 2 | 1 | 0 | 3 | 2 | 1 | 0 |
        // :---+---+---+---+---+---+---+---:
        // | 0 | x | x | x | 1 | x | x | x | T
        // | 0 | 0 | x | x | 0 | 1 | x | x | T
        // | 0 | 0 | 0 | x | 0 | 0 | 1 | x | T
        // | 0 | 0 | 0 | 0 | 0 | 0 | 0 | 1 | T
        // '---'---'---'---'---'---'---'---'            
        assign lt[i] =
            (~a[(i*4)+3] & ~a[(i*4)+2] & ~a[(i*4)+1] & ~a[(i*4)+0] & ~b[(i*4)+3] & ~b[(i*4)+2] & ~b[(i*4)+1] & b[(i*4)+0]) |
            (~a[(i*4)+3] & ~a[(i*4)+2] & ~a[(i*4)+1]               & ~b[(i*4)+3] & ~b[(i*4)+1] &  b[(i*4)+0]) |
            (~a[(i*4)+3] & ~a[(i*4)+2]                             & ~b[(i*4)+3] &  b[(i*4)+0]) |
            (~a[(i*4)+3]                                           &  b[(i*4)+3]);
        
        assign 
    
        end : LT_BLOCK
    endgenerate
    

    always @* begin
        casez({lt, gt, eq})
            {8'b1???_????, 8'b0???_????}: c = 1;
            {8'b01??_????, 8'b00??_????}: c = 1;
            {8'b001?_????, 8'b000?_????}: c = 1;
            {8'b0001_????, 8'b0000_????}: c = 1;
            {8'b0000_1???, 8'b0000_0???}: c = 1;
            {8'b0000_01??, 8'b0000_00??}: c = 1;
            {8'b0000_001?, 8'b0000_000?}: c = 1;
            {8'b0000_0001, 8'b0000_0000}: c = 1;
            default:                      c = 0;
        endcase
    end


endmodule : StructuralLogicalLT
`default_nettype wire