//------------------------------------------------------------------------
//
//
//------------------------------------------------------------------------
`default_nettype none
module Multiply
#(  //-----------------------------------//-------------------------------
    // Parameter(s)                      // Description(s)
    //-----------------------------------//-------------------------------
    parameter integer N         = 32,    // Data path width in bits
    parameter string  ALGORITHM = "RTL"  //
)  (//-----------------------------------//-------------------------------
    // Inputs                            // Description(s)
    //-----------------------------------//-------------------------------
    input wire [   N-1:0] a,             //
    input wire [   N-1:0] b,             //
    //-----------------------------------//-------------------------------
    // Outputs                           // Description(s)
    //-----------------------------------//-------------------------------
    output wire [2*N-1:0] c
);


    generate
        if (ALGORITHM == "RTL") begin
	     assign c = a * b;	
        end
    endgenerate
    

endmodule : Mutliply
`default_nettype wire

