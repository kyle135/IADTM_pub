//-----------------------------------------------------------------------------
// Licensing:   It's All Digital To Me (c) 2018 by Kyle D. Gilsdorf is licensed
//              under Creative Commons Attribution 4.0 International.
// Company:     It's All Digital To Me
// Engineer:    Kyle D. Gilsdorf (Kyle.Gilsdorf@asu.edu)
// IP Name:     FixedPointArithmetic
// Unit Name:   Add
// Algorithm:   PrefixAdd
// Modeling:    Behavioral
// Description: 
//-----------------------------------------------------------------------------
`default_nettype none
module BehavioralPrefixAdd
#(  //--------------------------//-----------------------------------------
    // Parameters               // Descriptions
    //--------------------------//-----------------------------------------
    parameter integer   N = 32  // Datapath width in bits
)  (//--------------------------//-----------------------------------------
    // Inputs                   // Descriptions
    //--------------------------//-----------------------------------------
    input  wire [N-1:0] a,      // Operand A
    input  wire [N-1:0] b,      // Operand B
    input  wire         ci,     // Carry in
    //--------------------------//-----------------------------------------
    // Outputs                  // Descriptions
    //--------------------------//-----------------------------------------
    output wire [N-1:0] c,      // Result
    output wire         co      // Carry out
);

//-------------------------------------------------------------------------
// Local Nets
//-------------------------------------------------------------------------

//-------------------------------------------------------------------------
// Continuous Assignments and Combinational Logic
//-------------------------------------------------------------------------

//-------------------------------------------------------------------------
// Synchronous Logic
//-------------------------------------------------------------------------

//-------------------------------------------------------------------------
// Module Instantiation
//-------------------------------------------------------------------------

endmodule : BehavioralPrefixAdd
`default_nettype wire
