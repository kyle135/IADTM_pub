`ifndef __BITWISESEQUENCER__SVH
    `define __BITWISESEQUENCER__SVH
//---------------------------------------------------------------------------------------
// Sequencer
//---------------------------------------------------------------------------------------
typedef uvm_sequencer #(BitWiseSequenceItem) BitWiseSequencer;
`endif // __BITWISESEQUENCER__SVH