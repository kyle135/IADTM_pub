`ifndef __UNARYSEQUENCER__SVH
    `define __UNARYSEQUENCER__SVH
//---------------------------------------------------------------------------------------
// Sequencer
//---------------------------------------------------------------------------------------
typedef uvm_sequencer #(UnarySequenceItem) UnarySequencer;
`endif // __UNARYSEQUENCER__SVH