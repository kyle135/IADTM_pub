

//-----------------------------------------------------------------------------
// SUM:
//     Truth Table                      K-Map
// .---.---.-----.---.  .------------.----------.---------.
// | a | b | cin | c |  |          c | cin' (0) | cin (1) |
// :---+---+-----+---:  :------------+----------+---------:
// | 0 | 0 |  0  | 0 |  | a' b' (00) |     0    |    1    | 
// | 0 | 0 |  1  | 1 |  :------------+----------+---------:   
// | 0 | 1 |  0  | 1 |  | a' b  (01) |     1    |    0    |  
// | 0 | 1 |  1  | 0 |  :------------+----------+---------:
// | 1 | 0 |  0  | 1 |  | a  b  (11) |     0    |    1    | 
// | 1 | 0 |  1  | 0 |  :------------+----------+---------:
// | 1 | 1 |  0  | 0 |  | a  b' (10) |     1    |    0    |
// | 1 | 1 |  1  | 1 |  '------------'----------'---------'
// '---'---'-----'---'
//
// SOP: c = (a'·b'·cin) + (a'·b·cin') + (a·b·cin) + (a·b'·cin') From the K-Map
//        = a·(b·cin + b'·cin') + a'·(b·cin' + b'·cin)
//        = a·~(B^C) + a'·(B^C)
//        = a ^ (b ^ c)
//        = a ^ b ^ c
//
//-----------------------------------------------------------------------------
// CARRY:
//     Truth Table                      K-Map
// .---.---.-----.------.  .------------.----------.---------.
// | a | b | cin | cout |  |       cout | cin' (0) | cin (1) |
// :---+---+-----+------:  :------------+----------+---------:
// | 0 | 0 |  0  |   0  |  | a' b' (00) |     0    |    0    | 
// | 0 | 0 |  1  |   0  |  :------------+----------+---------:   
// | 0 | 1 |  0  |   0  |  | a' b  (01) |     0    |    1    |  
// | 0 | 1 |  1  |   1  |  :------------+----------+---------:
// | 1 | 0 |  0  |   0  |  | a  b  (11) |     1    |    1    | 
// | 1 | 0 |  1  |   1  |  :------------+----------+---------:
// | 1 | 1 |  0  |   1  |  | a  b' (10) |     0    |    1    |
// | 1 | 1 |  1  |   1  |  '------------'----------'---------'
// '---'---'-----'------'
//
// SOP: cout = (b·cin) + (a·cin) + (a·b)
//           = cin·(a + b) + (a·b)
//-----------------------------------------------------------------------------
module RippleCarryAdder
#(  //--------------------------------------//---------------------------------
    // Parameters                           // Description(s)
    //--------------------------------------//---------------------------------
    parameter int    N     = 32,            // Datapath width in bits.
    parameter string MODEL = "Structural"   // Which modeling technique are we using?
)  (//--------------------------------------//---------------------------------
    // Inputs                               // Description(s)
    //--------------------------------------//---------------------------------
    input  wire [N-1:0] a,                  //
    input  wire [N-1:0] b,                  //
    input  wire         carry_in,           //
    //--------------------------------------//---------------------------------
    // Outputs                              // Description(s)
    //--------------------------------------//---------------------------------
    output wire [N-1:0] c,                  //
    output wire         carry_out           //
);
    
    //-------------------------------------------------------------------------
    // Local Signals
    //-------------------------------------------------------------------------

    //-------------------------------------------------------------------------
    // Combinational Logic
    //-------------------------------------------------------------------------
    
    //-------------------------------------------------------------------------
    // Sequential Logic
    //-------------------------------------------------------------------------

    //-------------------------------------------------------------------------
    // Module Instantiation
    //-------------------------------------------------------------------------
    generate
        if (MODEL == "Behavioral") begin : BEHAVIORAL_INTANSTIATION
            BehavioralRippleCarryAdder
            #(  //----------------------------------//---------------------------------
                // Parameters                       // Description(s)
                //----------------------------------//---------------------------------
                .N         ( N                   )  // Data-path width in bits
            )                                       //
            u_BehavioralRippleCarryAdder            //
            (   //----------------------------------//---------------------------------
                // Inputs                           // Direction, Size & Description(s)
                //----------------------------------//---------------------------------
                .a         ( a                   ), // [I][N] Operand A
                .b         ( b                   ), // [I][N] Operand B
                .carry_in  ( carry_in            ), // [I][1] Carry In
                //----------------------------------//---------------------------------
                // Outputs                          // Direction, Size & Description(s)
                //----------------------------------//---------------------------------
                .c         ( c                   ), // [O][N] Result Sum
                .carry_out ( carry_out           )  // [O][1] Result Carry
            );                                      //
        end : BEHAVIORAL_INTANSTIATION
        else if (MODEL == "DataFlow") begin : DATAFLOW_INTANSTIATION
            DataFlowRippleCarryAdder
            #(  //----------------------------------//---------------------------------
                // Parameters                       // Description(s)
                //----------------------------------//---------------------------------
                .N         ( N                   )  // Data-path width in bits
            )                                       //
            u_DataFlowRippleCarryAdder              //
            (   //----------------------------------//---------------------------------
                // Inputs                           // Direction, Size & Description(s)
                //----------------------------------//---------------------------------
                .a         ( a                   ), // [I][N] Operand A
                .b         ( b                   ), // [I][N] Operand B
                .carry_in  ( carry_in            ), // [I][1] Carry In
                //----------------------------------//---------------------------------
                // Outputs                          // Direction, Size & Description(s)
                //----------------------------------//---------------------------------
                .c         ( c                   ), // [O][N] Result Sum
                .carry_out ( carry_out           )  // [O][1] Result Carry
            );                                      //
        end : DATAFLOW_INTANSTIATION
        else if (MODEL == "Structural") begin : STRUCTURAL_INSTANTIATION
            StructuralRippleCarryAdder
            #(  //----------------------------------//---------------------------------
                // Parameters                       // Description(s)
                //----------------------------------//---------------------------------
                .N         ( N                   )  // Data-path width in bits
            )                                       //
            u_StructuralRippleCarryAdder            //
            (   //----------------------------------//---------------------------------
                // Inputs                           // Direction, Size & Description(s)
                //----------------------------------//---------------------------------
                .a         ( a                   ), // [I][N] Operand A
                .b         ( b                   ), // [I][N] Operand B
                .carry_in  ( carry_in            ), // [I][1] Carry In
                //----------------------------------//---------------------------------
                // Outputs                          // Direction, Size & Description(s)
                //----------------------------------//---------------------------------
                .c         ( c                   ), // [O][N] Result Sum
                .carry_out ( carry_out           )  // [O][1] Result Carry
            );                                      //
        end : STRUCTURAL_INSTANTIATION
    endgenerate

endmodule : RippleCarryAdder
