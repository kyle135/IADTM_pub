//---------------------------------------------------------------------------------------
// Licensing:       It's All Digital To Me © 2018 by Kyle D. Gilsdorf is licensed under
//                  Creative Commons Attribution 4.0 International 
//
// Company:         It's All Digital To Me
// Engineer:        Kyle D. Gilsdorf
// Module Name:     APB_hvl_pkg
// Description:
//---------------------------------------------------------------------------------------
package APB_hvl_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import APB_hdl_pkg::*;

    const logic FAILURE = 1'b0;
    const logic SUCCESS = 1'b1;

    `include "hvl/SequenceItems/src/APBSequenceItem.svh"
    `include "hvl/Config/src/APBConfig.svh"
    `include "hvl/Sequence/src/APBSequence.svh"
    `include "hvl/Sequencer/src/APBSequencer.svh"
    `include "hvl/Monitor/src/APBMonitor.svh"
    `include "hvl/Driver/src/APBDriver.svh"
    `include "hvl/Agent/src/APBAgent.svh"

endpackage : APB_hvl_pkg
