`ifndef __ADDSEQUENCER__SVH
    `define __ADDSEQUENCER__SVH
//---------------------------------------------------------------------------------------
// Sequencer
//---------------------------------------------------------------------------------------
typedef uvm_sequencer #(AddSequenceItem) AddSequencer;
`endif // __ADDSEQUENCER__SVH