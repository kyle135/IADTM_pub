


package ALU_hdl_pkg;


endpackage : ALU_hdl_pkg
