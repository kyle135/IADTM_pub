//---------------------------------------------------------------------------------------
// Company: It's All Digital To Me
// Engineer: Kyle D. Gilsdorf
// Create Date: 11/25/2020, 3:23:29 PM
//---------------------------------------------------------------------------------------
`default_nettype none
module StructuralCounter
#(  //------------------------------------------------------------------------------------
    //
    //------------------------------------------------------------------------------------

)  (//------------------------------------------------------------------------------------
    //
    //------------------------------------------------------------------------------------



);

endmodule : StructuralCounter
`default_nettype wire