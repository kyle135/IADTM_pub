



typedef enum logic [7:0] {
    R2000       = 1,
    R3000       = 2,
    R6000       = 3,
    R4000_R4400 = 4,

} Imp_t;


