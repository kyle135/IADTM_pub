//-----------------------------------------------------------------------------
// Licensing:    It's All Digital To Me © 2018 by Kyle D. Gilsdorf is licensed 
//               under Creative Commons Attribution 4.0 International.
// Company:      It's All Digital To Me
// Engineer:     Kyle D. Gilsdorf (Kyle.Gilsdorf@asu.edu)
//
//-----------------------------------------------------------------------------
`default_nettype none
module BehavioralCarrySaveAdd
#(  //--------------------------//---------------------------------------------
    // Parameters               // Description(s)
    //--------------------------//---------------------------------------------
    parameter integer   N = 32  //
)  (//--------------------------//---------------------------------------------
    // Inputs                   // Description(s)
    //--------------------------//---------------------------------------------
    input  wire [N-1:0] a,      //
    input  wire [N-1:0] b,      //
    input  wire         ci,     //
    //--------------------------//---------------------------------------------
    // Outputs                  // Description(s)
    //--------------------------//---------------------------------------------
    output reg  [N-1:0] c,      //
    output reg          co      //
);

    //-------------------------------------------------------------------------
    // Local Signals
    //-------------------------------------------------------------------------


    //-------------------------------------------------------------------------
    // Combinational Logic
    //-------------------------------------------------------------------------


endmodule : BehavioralCarrySaveAdd
`default_nettype wire
