`ifndef __LOGICALSEQUENCER__SVH
    `define __LOGICALSEQUENCER__SVH
//---------------------------------------------------------------------------------------
// Sequencer
//---------------------------------------------------------------------------------------
typedef uvm_sequencer #(LogicalSequenceItem) LogicalSequencer;
`endif // __LOGICALSEQUENCER__SVH