//---------------------------------------------------------------------------------------
// Company: It's All Digital To Me
// Engineer: Kyle D. Gilsdorf
// Create Date: 09/21/2013
// Design Name: Structural Logical Less Than (by n-bits)
// Unit Name: Logical
// Module Name: StructuralLogicalGT
// Project Name: BasicCombinationalLogic
// Dependencies: None
//
//  ¬x1 · y1 + 
// ¬(y1 ^ y1) ·  ¬x2 · y2 + 
// ¬(x1 ^ y1) · ¬(x2 ^ y2) ·  ¬x3 · y3
// ¬(x1 ^ y1) · ¬(x2 ^ y2) · ¬(x3 · y3) ·  ¬x4 · y4
//-----------------------------------------------------------------------------
`default_nettype none
module StructuralLogicalLT
#(  //----------------------------------//-------------------------------------
    // Parameter(s)                     // Description(s)
    //----------------------------------//-------------------------------------
    parameter integer N = 4             // The number of bits of the operands.
)  (//----------------------------------//-------------------------------------
    // Input(s)                         // Description(s)
    //----------------------------------//-------------------------------------
    input  wire [N-1:0] a,              // Operand A
    input  wire [N-1:0] b,              // Operand B
    //----------------------------------//-------------------------------------
    // Output(s)                        // Description(s)
    //----------------------------------//-------------------------------------
    output wire         c               // Result C
);

    //-------------------------------------------------------------------------
    // Local Signals
    //-------------------------------------------------------------------------
    wire [N-1:0] not_a;
    wire [N-1:0] not_a_and_b;
    wire [N-1:0] a_xor_b;
    wire [N-1:0] not_xor;
    wire [N-1:0] a_xor_b_and_chain;
    wire [N-1:0] a_xor_b_and_not_a_and_b_chain;
    wire [N-2:0] lt_chain;
    //-------------------------------------------------------------------------
    // Combinational Logic
    //-------------------------------------------------------------------------

    //-------------------------------------------------------------------------
    // Module instance(s)
    //-------------------------------------------------------------------------
    // a=0x9A48_810D ~a=0x65B7_7EF2
    // b=0x6222_8F65                                                        .
    //              .------.                                                |
    // a[31] -.----/|      |------------------------------------------------|
    //        |     | ¬a·b |                                                |
    // b[31] -|--.--|      |                                                |
    //        |  |  '------'.-----.                                         |
    //        |  '----------|     |-.                                       |
    //        |             | a^b | |                                       |
    //        '-------------|     | |  .------.                             |
    //                      '-----' '-/|      |-----------------------------|
    //           .------.              | ¬a·b |
    //   a[30] -/|      |--------------|      |
    //           | ¬a·b |              '------'
    //   b[30] --|      |
    //           '------'

    //           .------.
    //   a[30] -/|      |
    //           | ¬a·b |
    //   b[30] --|      |
    //           '------'  
    //                   
    //
    // (a < b ) =                                                          (~a[31] · b[31])  + 
    //           (~(a[31] ^ b[31])                                       & (~a[30] · b[30])) + 
    //           (~(a[31] ^ b[31]) & ~(a[30] ^ b[30])                    & (~a[29] · b[29])) +
    //           (~(a[31] ^ b[31]) & ~(a[30] ^ b[30]) & ~(a[30] ^ b[30]) & (~a[28] · b[28])) +
    // .----.------.-------.------.--------------.-------------.----------------.
    // |  i | a[i] | ~a[i] | b[i] | ~a[i] · b[i] | a[i] ^ b[i] | ~(a[i] ^ b[i]) | a[i] < b[i] |
    // :----+------+-------+------'--------------+-------------+----------------+-------------:
    // | 15 |  1   |   0   |  1   |       0      |      0      |        1       | 0 +
    // | 14 |  0   |   1   |  0   |       0      |      0      |        1       | 0     0
    // | 13 |  0   |   1   |  1   |       1      |      1      |        0       |      0
    // | 12 |  0   |   1   |  0   |       0      |      0      |        1       |      0
    // | 11 |  0   |   1   |  0   |       0      |      0      |        1       |      0
    // | 10 |  0   |   1   |  1   |       1      |      1      |        0       |      0
    // |  9 |  0   |   1   |  1   |       1      |      1      |        0       |      0
    // |  8 |  1   |   0   |  0   |       0      |      1      |        0       |      0
    // |  7 |  0   |   1   |  1   |       1      |      1      |        0       |      
    // |  7 |  0   |   1   |  1   |       1      |      1      |        0       |
    // |  6 |  0   |   1   |  1   |       1      |      1      |        0       |
    // |  5 |  0   |   1   |  1   |       1      |      1      |        0       |    0
    // |  4 |  0   |   1   |  0   |       0      |      0      |        1       |    0
    // |  3 |  1   |   0   |  0   |       0      |      1      |        0       |    0
    // |  2 |  1   |   0   |  0   |       0      |      1      |        0       |    0
    // |  1 |  0   |   1   |  1   |       1      |      1      |        0       |    0
    // |  0 |  1   |   0   |  1   |       0      |      0      |        1       |    0    
    // '----'------'-------'------'--------------'-------------'----------------'

    genvar i;
    generate
        for (i = N-1; i >= 0 ; i = i - 1) begin : LT_BLOCK
            //  ¬x1 · y1 + 
            // \___/
            not u_not_a (not_a[i], a[i]);
            //  ¬x1 · y1 + 
            // \________/
            and u_not_a_and_b (not_a_and_b[i], not_a[i], b[i]);
            // ¬(x1 ^ y1) · ¬(x2 ^ y2) · ¬(x3 · y3) ...
            //  \_______/    \_______/    \_______/
            xor u_a_xor_b (a_xor_b[i], a[i], b[i]);
            // ¬(x1 ^ y1) · ¬(x2 ^ y2) · ¬(x3 · y3) ...
            //\__________/ \__________/ \__________/
            not u_not_xor (not_xor[i], a_xor_b[i]);
            // i = 0   ...
            // i = 1   ¬(y1 ^ y1) ·  ...
            //        \__________/
            // i = 2   ¬(x1 ^ y1) · ¬(x2 ^ y2) · ...
            //        \__________/ \__________/
            // i = 3   ¬(x1 ^ y1) · ¬(x2 ^ y2) · ¬(x3 ^ y3) · ...
            //        \__________/ \__________/ \__________/
            and u_not_a_xor_b_and_chain(a_xor_b_and_chain[i], not_xor[i], a_xor_b_and_chain[N-1:i+1]);

            and u_a_xor_b_and_not_a_and_b_chain(
                a_xor_b_and_not_a_and_b_chain[i], 
                a_xor_b_and_chain[i],
                not_a_and_b[i]);


            if (i == N-1) begin
                or u_or_lt_chain(c, lt_chain[i+1], a_xor_b_and_not_a_and_b_chain[i]);
            end else begin
                or u_or_lt_chain(lt_chain[i], lt_chain[i+1], a_xor_b_and_not_a_and_b_chain[i]);
            end
        end : LT_BLOCK
    endgenerate

endmodule : StructuralLogicalLT
`default_nettype wire