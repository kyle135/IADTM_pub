module FixedPointDivide
#(  //-------------------------------------------
    //
    //--------------------------------
    parameter integer N = 32
)  (//--------------------------------
    //
    //-----------------------------------------
    input  wire [N-1:0] a,
	input  wire [N-1:0] b,
    //-----------------------------------------
    //
    //-----------------------------------------
	output wire [2*N-1:0] c
);


    assign c = a / b;


endmodule : FixedPointDivide
