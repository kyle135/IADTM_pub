


`default_nettype none
module DataFlowLogicalOR
#(  //----------------------------------//-------------------------------------
    // Parameters                       // Description(s)
    //----------------------------------//-------------------------------------    
    parameter integer N = 8             // Width of operands and result in bits
)  (//----------------------------------//-------------------------------------
    // Input Ports                      // Description(s)
    //----------------------------------//-------------------------------------
    input  wire [N-1:0] a,              // Operand A
    input  wire [N-1:0] b,              // Operand B
    //----------------------------------//-------------------------------------    
    // Output Ports                     // Description(s)
    //----------------------------------//-------------------------------------
    output wire            c            // Result C
);
    //----------------------------------//-------------------------------------
    // Local Signals                    // Description(s)
    //----------------------------------//-------------------------------------
    wire [N-1:0] a_or;                  //
    wire [N-1:0] b_or;                  //
    
    
    //----------------------------------//-------------------------------------
    // Combinational Logic              // Description(s)
    //----------------------------------//-------------------------------------    
    assign a_or = |a;
    assign b_or = |b;
    assign c    = a_or | b_or;


endmodule : DataFlowLogicalOR
`default_nettype wire
